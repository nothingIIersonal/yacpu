﻿`ifndef HWID_VH
`define HWID_VH


parameter HWID_SCNP                  = 2'b00;
parameter HWID_CPU                   = 2'b01;
parameter HWID_GPU                   = 2'b10;
parameter HWID_PERIPHERAL_CONTROLLER = 2'b11;


`endif