/*
 * Copyright (C) 2022 nothingIIersonal.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */



`timescale 1ns / 1ps



/*
 *   __     __      __  __  _____ _    _ 
 *   \ \   / //\   |  \/  |/ ____| |  | |
 *    \ \_/ //  \  | \  / | |    | |  | |
 *     \   // /\ \ | |\/| | |    | |  | |
 *      | |/ ____ \| |  | | |____| |__| |
 *      |_/_/    \_\_|  |_|\_____|\____/
 *
 *
 * UART TX module
 *
 * Designer : Magomedov R. M. (https://github.com/nothingIIersonal)
 * Designer : Glazunov  N. M. (https://github.com/nikikust        )
 *
 */



module uart_tx
#
(
    parameter CLK_RATE_MHz      =   100,
    parameter DATA_WIDTH        =     8,
    parameter CLK_COUNTER_WIDTH =    14,
    parameter COUNTER_REG_WIDTH =     4,
    parameter CLK_COUNTER_INV   = 10416,
    parameter BOUDRATE          =  9600
)
(
    input  wire                        clk_in,
    input  wire                        rst_in,

    input  wire                        tx_en_in,

    input  wire [DATA_WIDTH - 1: 0]    txdata_in,

    output reg                         tx_out,
    output reg                         done_transmit_out
);

    reg                            state_reg;

    reg [COUNTER_REG_WIDTH: 0]     counter_reg;
    reg [CLK_COUNTER_WIDTH: 0]     clk_counter;

    reg                            tx_en_in_reg;
    reg                            tx_en_in_flag_reg;

    reg [DATA_WIDTH - 1: 0]        txdata_in_reg;

    reg                            clk_tx;


    localparam // state_regs
        START_TRANSMIT = 1'h0,
        SEND_DATA      = 1'h1;


    initial
    begin
        state_reg         <= START_TRANSMIT;

        counter_reg       <= {COUNTER_REG_WIDTH + 1'b1{1'b0}};
        clk_counter       <= {CLK_COUNTER_WIDTH + 1'b1{1'b0}};

        tx_en_in_reg      <= 1'b0;
        tx_en_in_flag_reg <= 1'b0;

        txdata_in_reg     <= {DATA_WIDTH{1'b1}};

        clk_tx            <= 1'b0;

        tx_out            <= 1'b1;

        done_transmit_out <= 1'b1;
    end


    always @(posedge clk_in)
    begin
        ////
        // Process enable and stop transmission signals
        if (tx_en_in && done_transmit_out) begin
            tx_en_in_reg      <= 1'b1;
            txdata_in_reg     <= txdata_in;
            done_transmit_out <= 1'b0;
        end else if (tx_en_in_flag_reg) begin
            tx_en_in_reg      <= 1'b0;
        end
        ////


        if (!rst_in) begin
            ////
            // Generate TX clock
            if (clk_counter < CLK_COUNTER_INV) begin
                clk_tx      <= 1'b0;
                clk_counter <= clk_counter + {{CLK_COUNTER_WIDTH{1'b0}}, 1'b1};
            end else begin
                clk_counter <= {CLK_COUNTER_WIDTH + 1'b1{1'b0}};
                clk_tx      <= 1'b1;
            end
            ////

            ////
            // Send data process
            if (clk_tx) begin
                case (state_reg)
                    START_TRANSMIT: begin
                        if (tx_en_in_reg) begin                
                            state_reg         <= SEND_DATA;
                            tx_en_in_flag_reg <= 1'b1;
                            tx_out            <= 1'b0;
                        end
                    end
                    SEND_DATA: begin
                        tx_en_in_flag_reg     <= 1'b0;

                        if (counter_reg <= DATA_WIDTH - 1) begin
                            tx_out            <= txdata_in_reg[counter_reg[COUNTER_REG_WIDTH - 1: 0]];
                            counter_reg       <= counter_reg + {{COUNTER_REG_WIDTH{1'b0}}, 1'b1};
                        end else begin
                            state_reg         <= START_TRANSMIT;

                            txdata_in_reg     <= {DATA_WIDTH{1'b1}};
                            tx_out            <= 1'b1;
                            counter_reg       <= {COUNTER_REG_WIDTH + 1'b1{1'b0}};
                            done_transmit_out <= 1'b1;
                        end
                    end
                endcase
            end
            /////
        end else begin
            state_reg         <= START_TRANSMIT;

            counter_reg       <= {COUNTER_REG_WIDTH + 1'b1{1'b0}};
            clk_counter       <= {CLK_COUNTER_WIDTH + 1'b1{1'b0}};

            txdata_in_reg     <= {DATA_WIDTH{1'b1}};

            clk_tx            <= 1'b0;

            tx_out            <= 1'b1;

            done_transmit_out <= 1'b1;
        end
    end

endmodule
