﻿`timescale 1ns / 1ps


module uart_tx
(
    input  wire in_clk
)


endmodule
