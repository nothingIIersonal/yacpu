`ifndef PARAMETERS_VH
`define PARAMETERS_VH


// `define DEBUG


// GLOBAL
parameter SYSTEM_CLOCK_MHz  =   100;
parameter UART_BAUDRATE     = 57600;
//// GLOBAL


// MEMORY
parameter MEMORY_WORD_WIDTH =    8;
parameter MEMORY_CAPACITY   = 1024;
//// MEMORY


`endif
